Library IEEE;
USE ieee.std_logic_1164.all;
USE ieee.numeric_std.all;

PACKAGE ADF IS
	TYPE TAB IS ARRAY (NATURAL RANGE <>) OF INTEGER; -- tableau de integer
END PACKAGE;
